`include "defines.v"

module openmips(

	input	wire										clk,
	input wire										rst,
	
 
	input wire[`RegBus]           rom_data_i,
	output wire[`RegBus]           rom_addr_o,
	output wire                    rom_ce_o,

	//连接data_ram
	input wire[`RegBus]           ram_data_i,
	output wire[`RegBus]           ram_addr_o,
	output wire[`RegBus]           ram_data_o,
	output wire                    ram_we_o,
	output wire[3:0]               ram_sel_o,
	output wire[3:0]               ram_ce_o
	
);

	// 参数定义说明
	// xx_o----->某一个模块的输出,如ex_wd_o表示ex模块的输出
	// xx_i----->某一个模块的输入,如ex_wd_o表示ex模块的输入


    //IF/ID模块与译码阶段ID模块
	wire[`InstAddrBus] pc;
	wire[`InstAddrBus] id_pc_i;
	wire[`InstBus] id_inst_i;
	
	//连接译码阶段ID模块的输出与ID/EX模块的输入
	wire[`AluOpBus] id_aluop_o;
	wire[`AluSelBus] id_alusel_o;
	wire[`RegBus] id_reg1_o;
	wire[`RegBus] id_reg2_o;
	wire id_wreg_o;
	wire[`RegAddrBus] id_wd_o;
	
	//连接ID/EX模块的输出与执行阶段EX模块的输入
	wire[`AluOpBus] ex_aluop_i;
	wire[`AluSelBus] ex_alusel_i;
	wire[`RegBus] ex_reg1_i;
	wire[`RegBus] ex_reg2_i;
	wire ex_wreg_i;
	wire[`RegAddrBus] ex_wd_i;
	
	//连接执行阶段EX模块的输出与EX/MEM模块的输入
	wire ex_wreg_o;
	wire[`RegAddrBus] ex_wd_o;
	wire[`RegBus] ex_wdata_o;
	//Hilo
	wire ex_whilo_o;
	wire[`RegBus] ex_hi_o;
	wire[`RegBus] ex_lo_o;


	//连接EX/MEM模块的输出与访存阶段MEM模块的输入
	wire mem_wreg_i;
	wire[`RegAddrBus] mem_wd_i;
	wire[`RegBus] mem_wdata_i;
	//Hilo
	wire mem_whilo_i;
	wire[`RegBus] mem_hi_i;
	wire[`RegBus] mem_lo_i;

	//连接访存阶段MEM模块的输出与MEM/WB模块的输入
	wire mem_wreg_o;
	wire[`RegAddrBus] mem_wd_o;
	wire[`RegBus] mem_wdata_o;
	//Hilo
	wire mem_whilo_o;
	wire[`RegBus] mem_hi_o;
	wire[`RegBus] mem_lo_o;

	
	//连接MEM/WB模块的输出与回写阶段的输入	
	wire wb_wreg_i;
	wire[`RegAddrBus] wb_wd_i;
	wire[`RegBus] wb_wdata_i;
	//连接MEM/WB模块与Hilo
	wire hilo_we_i;
	wire[`RegBus] hi_i;
	wire[`RegBus] lo_i;
	
	//连接译码阶段ID模块与通用寄存器Regfile模块
	wire reg1_read;
	wire reg2_read;
	wire[`RegBus] reg1_data;
	wire[`RegBus] reg2_data;
	wire[`RegAddrBus] reg1_addr;
	wire[`RegAddrBus] reg2_addr;

	//连接回写阶段HELO与执行阶段
	wire[`RegBus] hi_o;
	wire[`RegBus] lo_o;

	// ctrl 
	wire[5:0] stall;
	wire      stallreq_from_id_i;
	wire      stallreq_from_ex_i;

	//div
	wire[`DoubleRegBus] div_result_i; // 64位
	wire          div_ready_i;
	wire          signed_div_i;
	wire[`RegBus] div_opdata1_i;
	wire[`RegBus] div_opdata2_i;
	wire          div_start_i;

	// 分支跳转
	wire branch_flag;
	wire[`InstAddrBus]    branch_target_address;
	wire                  id_is_in_delayslot;  //这条在译码的时候发现为延迟槽指令，is_in_delayslot为true
	wire                  next_inst_in_delayslot; // 现在处于译码的指令是分支跳转指令并且满足跳转条件     
	wire[`RegBus]         id_link_address;  // 需要保存的返回地址
	wire                  id_ex_is_in_delayslot;
	wire[`RegBus]         ex_link_address;
	wire                  ex_is_in_delayslot;  // 这个暂时没有用
  
  //pc_reg例化
	pc_reg pc_reg0(
		.clk(clk),
		.rst(rst),

		// 分支跳转指令增加的接口
		.branch_flag_i(branch_flag),
		.branch_target_address_i(branch_target_address),

		.pc(pc),
		.stall(stall),
		.ce(rom_ce_o)	
	);
	
  assign rom_addr_o = pc;

  //通用寄存器Regfile例化
	regfile regfile1(
		.clk (clk),
		.rst (rst),
		.we	(wb_wreg_i),  // 是否要写,最终信号传入寄存器堆
		.waddr (wb_wd_i),
		.wdata (wb_wdata_i),
		.re1 (reg1_read),
		.raddr1 (reg1_addr),
		.rdata1 (reg1_data),
		.re2 (reg2_read),
		.raddr2 (reg2_addr),
		.rdata2 (reg2_data)
	);

	hilo_reg hilo_reg0(
		.clk(clk),
		.rst(rst),
		// 写
		.we(hilo_we_i),
		.hi_i(hi_i),
		.lo_i(lo_i),
		// 读
        .hi_o(hi_o),
        .lo_o(lo_o)
	);

	// div模块
	div div0(
		.clk(clk),
		.rst(rst),
	
		.signed_div_i(signed_div_i),
		.opdata1_i(div_opdata1_i),
		.opdata2_i(div_opdata2_i),
		.start_i(div_start_i),
		.annul_i(1'b0),
	
		.result_o(div_result_i),
		.ready_o(div_ready_i)
	);

	ctrl ctrl0(
		.rst(rst),
		.stallreq_from_id(stallreq_from_id_i),
		.stallreq_from_ex(stallreq_from_ex_i),
		.stall(stall)       	
	);

  //IF/ID模块例化
	if_id if_id0(
		.clk(clk),
		.rst(rst),
		.if_pc(pc),
		.stall(stall),
		.if_inst(rom_data_i),
		.id_pc(id_pc_i),
		.id_inst(id_inst_i)      	
	);
	
	//译码阶段ID模块
	id id0(
		.rst(rst),
		.pc_i(id_pc_i),
		.inst_i(id_inst_i),

		.stallreq(stallreq_from_id_i),

		// 分支跳转指令增加的接口
		.is_in_delayslot_i(id_is_in_delayslot),  //这条在译码的时候发现为延迟槽指令，is_in_delayslot为true
		.next_inst_in_delayslot_o(next_inst_in_delayslot), // 现在处于译码的指令是分支跳转指令并且满足跳转条件
		.branch_flag_o(branch_flag),
		.branch_target_address_o(branch_target_address),       
		.link_addr_o(id_link_address),  // 需要保存的返回地址
		.is_in_delayslot_o(id_ex_is_in_delayslot),

		//处于执行阶段的指令要写入的目的寄存器信息
		.ex_wreg_i(ex_wreg_o),
		.ex_wdata_i(ex_wdata_o),
		.ex_wd_i(ex_wd_o),
	
		//处于访存阶段的指令要写入的目的寄存器信息
		.mem_wreg_i(mem_wreg_o),
		.mem_wdata_i(mem_wdata_o),
		.mem_wd_i(mem_wd_o),

		.reg1_data_i(reg1_data),
		.reg2_data_i(reg2_data),

		//送到regfile的信息
		.reg1_read_o(reg1_read),
		.reg2_read_o(reg2_read), 	  

		.reg1_addr_o(reg1_addr),
		.reg2_addr_o(reg2_addr), 
	  	
		//送到ID/EX模块的信息
		.aluop_o(id_aluop_o),
		.alusel_o(id_alusel_o),
		.reg1_o(id_reg1_o),
		.reg2_o(id_reg2_o),
		.wd_o(id_wd_o),
		.wreg_o(id_wreg_o)
	);

	

	//ID/EX模块
	id_ex id_ex0(
		.clk(clk),
		.rst(rst),

		.id_link_address(id_link_address),
		.id_is_in_delayslot(id_is_in_delayslot),
		.next_inst_in_delayslot_i(next_inst_in_delayslot),	
		.ex_link_address(ex_link_address),
		.ex_is_in_delayslot(ex_is_in_delayslot),
		.is_in_delayslot_o(id_ex_is_in_delayslot),
		
		
		//从译码阶段ID模块传递的信息
		.id_aluop(id_aluop_o),
		.id_alusel(id_alusel_o),
		.id_reg1(id_reg1_o),
		.id_reg2(id_reg2_o),
		.id_wd(id_wd_o),
		.id_wreg(id_wreg_o),

		.stall(stall),
	
		//传递到执行阶段EX模块的信息
		.ex_aluop(ex_aluop_i),
		.ex_alusel(ex_alusel_i),
		.ex_reg1(ex_reg1_i),
		.ex_reg2(ex_reg2_i),
		.ex_wd(ex_wd_i),
		.ex_wreg(ex_wreg_i)
	);		
	
	//EX模块
	ex ex0(
		.rst(rst),

		//送到执行阶段EX模块的信息
		.aluop_i(ex_aluop_i),
		.alusel_i(ex_alusel_i),
		.reg1_i(ex_reg1_i),
		.reg2_i(ex_reg2_i),
		.wd_i(ex_wd_i),
		.wreg_i(ex_wreg_i),

		//是否转移、以及link address
		.link_address_i(ex_link_address),
		.is_in_delayslot_i(ex_is_in_delayslot),  // 这个暂时没有用

		// 因为数据移动指令(HILO)而添加的接口
		.hi_i(hi_o),  // 对应Hilo寄存器的值
		.lo_i(lo_o),
		.mem_whilo_i(mem_whilo_o),  // 处于访存阶段的指令是不是要写Hilo
		.mem_hi_i(mem_hi_o),  // 访存阶段要写入hi寄存器的值
		.mem_lo_i(mem_lo_o),  // 访存阶段要写入lo寄存器的值
		.wb_whilo_i(hilo_we_i),  // 处于写回阶段的指令是不是要写Hilo
		.wb_hi_i(hi_i),  // 写回阶段要写入hi寄存器的值
		.wb_lo_i(lo_i),  // 写回阶段要写入lo寄存器的值
		.whilo_o(ex_whilo_o),  // 是否要写Hilo
		.hi_o(ex_hi_o),  // 写入hi的值 
		.lo_o(ex_lo_o),  // 写入lo的值

		//div
		.div_result_i(div_result_i),
		.div_ready_i(div_ready_i),
		.stallreq(stallreq_from_ex_i),
		.div_opdata1_o(div_opdata1_i),
		.div_opdata2_o(div_opdata2_i),
		.div_start_o(div_start_i),
		.signed_div_o(signed_div_i),

	  	//EX模块的输出到EX/MEM模块信息
		.wd_o(ex_wd_o),
		.wreg_o(ex_wreg_o),
		.wdata_o(ex_wdata_o)
		
	);

  //EX/MEM模块
  ex_mem ex_mem0(
		.clk(clk),
		.rst(rst),
	  
		//来自执行阶段EX模块的信息	
		.ex_wd(ex_wd_o),
		.ex_wreg(ex_wreg_o),
		.ex_wdata(ex_wdata_o),

		.stall(stall),
	
		// Hilo寄存器添加的接口
		.ex_whilo(ex_whilo_o),
		.ex_hi(ex_hi_o),
		.ex_lo(ex_lo_o),
		.mem_whilo(mem_whilo_i),
		.mem_hi(mem_hi_i),
		.mem_lo(mem_lo_i),

		//送到访存阶段MEM模块的信息
		.mem_wd(mem_wd_i),
		.mem_wreg(mem_wreg_i),
		.mem_wdata(mem_wdata_i)

						       	
	);
	
  //MEM模块例化
	mem mem0(
		.rst(rst),
	
		//来自EX/MEM模块的信息	
		.wd_i(mem_wd_i),
		.wreg_i(mem_wreg_i),
		.wdata_i(mem_wdata_i),

		// Hilo寄存器添加的接口
		.whilo_i(mem_whilo_i),
		.hi_i(mem_hi_i),
		.lo_i(mem_lo_i),
		.whilo_o(mem_whilo_o),
		.hi_o(mem_hi_o),
		.lo_o(mem_lo_o),
	  
		//送到MEM/WB模块的信息
		.wd_o(mem_wd_o),
		.wreg_o(mem_wreg_o),
		.wdata_o(mem_wdata_o),

		//memory与mem相连
		.mem_data_i(ram_data_i),
		.mem_addr_o(ram_addr_o),
		.mem_we_o(ram_we_o),
		.mem_sel_o(ram_sel_o),
		.mem_data_o(ram_data_o),
		.mem_ce_o(ram_ce_o)
	);

  //MEM/WB模块
	mem_wb mem_wb0(
		.clk(clk),
		.rst(rst),

		//来自访存阶段MEM模块的信息	
		.mem_wd(mem_wd_o),
		.mem_wreg(mem_wreg_o),
		.mem_wdata(mem_wdata_o),

		.stall(stall),

		// Hilo寄存器添加的接口
		.mem_whilo(mem_whilo_o),
		.mem_hi(mem_hi_o),
		.mem_lo(mem_lo_o),
		.wb_whilo(hilo_we_i),
		.wb_hi(hi_i),
		.wb_lo(lo_i),
		
		//送到回写阶段的信息
		.wb_wd(wb_wd_i),
		.wb_wreg(wb_wreg_i),
		.wb_wdata(wb_wdata_i)
									       	
	);

endmodule